[0m[[0m[0minfo[0m] [0m[0mwelcome to sbt 1.10.2 (N/A Java 23.0.1-internal)[0m[0J
[0J[0m[[0m[0minfo[0m] [0m[0mloading settings for project chisel-build from plugins.sbt ...[0m[0J
[0J[0m[[0m[0minfo[0m] [0m[0mloading project definition from /users/students/r0886198/snax_cluster/hw/chisel/project[0m[0J
[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[1000D
[2K[2K  | => chisel-build / dependencyPositions 0s
[2K[2A[1000D[0J[0J[0J[1000D
[2K[2K  | => chisel-build / Compile / compileIncremental 0s
[2K[2A[1000D[0J[0m[[0m[0minfo[0m] [0m[0mloading settings for project root from build.sbt ...[0m[0J
[0J[0m[[0m[0minfo[0m] [0m[0mset current project to snax-streamer (in build file:/users/students/r0886198/snax_cluster/hw/chisel/)[0m[0J
[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[0J[1000D
[2K[2K  | => root / scalaCompilerBridgeBinaryJar 0s
[2K  | => root / update 0s
[2K[3A[1000D[1000D
[2K
[2K[2K  | => root / scalaCompilerBridgeBinaryJar 0s
[2K[3A[1000D[1000D
[2K
[2K[2K  | => root / scalaCompilerBridgeBinaryJar 0s
[2K[3A[1000D[1000D
[2K
[2K[2K  | => root / scalaCompilerBridgeBinaryJar 0s
[2K[3A[1000D[1000D
[2K
[2K[2K  | => root / scalaCompilerBridgeBinaryJar 0s
[2K[3A[1000D[0m[[0m[0minfo[0m] [0m[0mcompiling 2 Scala sources to /users/students/r0886198/snax_cluster/hw/chisel/target/scala-2.13/classes ...[0m[0J
[0J[1000D
[2K[2K  | => root / scalaCompilerBridgeBinaryJar 0s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / compileIncremental 0s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / compileIncremental 1s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / compileIncremental 2s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / compileIncremental 3s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / compileIncremental 4s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / compileIncremental 5s
[2K[2A[1000D[0J[1000D
[2K[2K  | => root / Compile / packageBin 0s
[2K[2A[1000D[1000D
[2K[2K  | => root / Compile / bgRunMain 0s
[2K[2A[1000D[0J[0m[[0m[0minfo[0m] [0m[0mrunning snax.DataPathExtension.RescaleDownEmitter [0m[0J
[0J[[33mwarn[0m] src/main/scala/snax/DataPathExtension/RescaleDown.scala 141:13: [W004] Dynamic index with width 7 is too wide for Vec of size 48 (expected index width 6).[0J
[[33mwarn[0m]         regs(counter.io.value * (extensionParam.dataWidth / in_elementWidth).U + i.U) := PE.io.data_o.asSInt[0J
[[33mwarn[0m]             ^[0J
[0J[[33mwarn[0m] There were [33m1 warning(s)[0m during hardware elaboration.[0J
[0J// Generated by CIRCT firtool-1.62.0[0J
// Standard header to adapt well known macros for register randomization.[0J
`ifndef RANDOMIZE[0J
  `ifdef RANDOMIZE_REG_INIT[0J
    `define RANDOMIZE[0J
  `endif // RANDOMIZE_REG_INIT[0J
`endif // not def RANDOMIZE[0J
[0J
// RANDOM may be set to an expression that produces a 32-bit random unsigned value.[0J
`ifndef RANDOM[0J
  `define RANDOM $random[0J
`endif // not def RANDOM[0J
[0J
// Users can define INIT_RANDOM as general code that gets injected into the[0J
// initializer block for modules with registers.[0J
`ifndef INIT_RANDOM[0J
  `define INIT_RANDOM[0J
`endif // not def INIT_RANDOM[0J
[0J
// If using random initialization, you can also define RANDOMIZE_DELAY to[0J
// customize the delay used, otherwise 0.002 is used.[0J
`ifndef RANDOMIZE_DELAY[0J
  `define RANDOMIZE_DELAY 0.002[0J
`endif // not def RANDOMIZE_DELAY[0J
[0J
// Define INIT_RANDOM_PROLOG_ for use in our modules below.[0J
`ifndef INIT_RANDOM_PROLOG_[0J
  `ifdef RANDOMIZE[0J
    `ifdef VERILATOR[0J
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM[0J
    `else  // VERILATOR[0J
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end[0J
    `endif // VERILATOR[0J
  `else  // RANDOMIZE[0J
    `define INIT_RANDOM_PROLOG_[0J
  `endif // RANDOMIZE[0J
`endif // not def INIT_RANDOM_PROLOG_[0J
[0J
// Include register initializers in init blocks unless synthesis is set[0J
`ifndef SYNTHESIS[0J
  `ifndef ENABLE_INITIAL_REG_[0J
    `define ENABLE_INITIAL_REG_[0J
  `endif // not def ENABLE_INITIAL_REG_[0J
`endif // not def SYNTHESIS[0J
[0J
// Include rmemory initializers in init blocks unless synthesis is set[0J
`ifndef SYNTHESIS[0J
  `ifndef ENABLE_INITIAL_MEM_[0J
    `define ENABLE_INITIAL_MEM_[0J
  `endif // not def ENABLE_INITIAL_MEM_[0J
`endif // not def SYNTHESIS[0J
[0J
module DataPathExtension_Demux_W512(	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:45[0J
  output         io_in_ready,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  input          io_in_valid,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  input  [511:0] io_in_bits,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  input          io_out_0_ready,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  output         io_out_0_valid,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  output [511:0] io_out_0_bits,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  input          io_out_1_ready,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  output         io_out_1_valid,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  output [511:0] io_out_1_bits,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
  input          io_sel	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:9:14[0J
);[0J
[0J
  assign io_in_ready = io_sel ? io_out_1_ready : ~io_sel & io_out_0_ready;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:45, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:15:15, :19:{17,26}, :21:23[0J
  assign io_out_0_valid = ~io_sel & io_in_valid;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:45, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:19:{17,26}, :20:23, :23:23[0J
  assign io_out_0_bits = io_in_bits;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:45[0J
  assign io_out_1_valid = io_sel & io_in_valid;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:45, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:19:26, :20:23, :23:23[0J
  assign io_out_1_bits = io_in_bits;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:45[0J
endmodule[0J
[0J
module DataPathExtension_Mux_W512(	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:44[0J
  output         io_in_0_ready,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  input          io_in_0_valid,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  input  [511:0] io_in_0_bits,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  output         io_in_1_ready,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  input          io_in_1_valid,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  input  [511:0] io_in_1_bits,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  input          io_out_ready,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  output         io_out_valid,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  output [511:0] io_out_bits,	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
  input          io_sel	// src/main/scala/snax/utils/MuxDemuxDecoupled.scala:89:14[0J
);[0J
[0J
  assign io_in_0_ready = ~io_sel & io_out_ready;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:44, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:99:{17,26}, :101:22, :104:22[0J
  assign io_in_1_ready = io_sel & io_out_ready;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:44, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:99:26, :101:22, :104:22[0J
  assign io_out_valid = io_sel ? io_in_1_valid : ~io_sel & io_in_0_valid;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:44, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:95:16, :99:{17,26}, :100:22[0J
  assign io_out_bits = io_sel ? io_in_1_bits : io_in_0_bits;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:44, src/main/scala/snax/utils/MuxDemuxDecoupled.scala:99:26, :102:22[0J
endmodule[0J
[0J
module RescaleDownCounter(	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
  input        clock,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
               reset,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
               io_tick,	// src/main/scala/snax/utils/Counter.scala:14:21[0J
               io_reset,	// src/main/scala/snax/utils/Counter.scala:14:21[0J
  output [1:0] io_value	// src/main/scala/snax/utils/Counter.scala:14:21[0J
);[0J
[0J
  reg [1:0] value;	// src/main/scala/snax/utils/Counter.scala:24:26[0J
  always @(posedge clock or posedge reset) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
    if (reset)	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
      value <= 2'h0;	// src/main/scala/snax/utils/Counter.scala:24:26, :30:25[0J
    else if (io_reset)	// src/main/scala/snax/utils/Counter.scala:14:21[0J
      value <= 2'h0;	// src/main/scala/snax/utils/Counter.scala:24:26, :30:25[0J
    else if (io_tick) begin	// src/main/scala/snax/utils/Counter.scala:14:21[0J
      if (value != 2'h3)	// src/main/scala/snax/utils/Counter.scala:24:26, :30:{32,42}, :39:38[0J
        value <= value + 2'h1;	// src/main/scala/snax/utils/Counter.scala:24:26, :30:55[0J
      else	// src/main/scala/snax/utils/Counter.scala:30:32[0J
        value <= 2'h0;	// src/main/scala/snax/utils/Counter.scala:24:26, :30:25[0J
    end[0J
  end // always @(posedge, posedge)[0J
  `ifdef ENABLE_INITIAL_REG_	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
    `ifdef FIRRTL_BEFORE_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
      `FIRRTL_BEFORE_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
    `endif // FIRRTL_BEFORE_INITIAL[0J
    initial begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
      automatic logic [31:0] _RANDOM[0:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
      `ifdef INIT_RANDOM_PROLOG_	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
        `INIT_RANDOM_PROLOG_	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
      `endif // INIT_RANDOM_PROLOG_[0J
      `ifdef RANDOMIZE_REG_INIT	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
        _RANDOM[/*Zero width*/ 1'b0] = `RANDOM;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
        value = _RANDOM[/*Zero width*/ 1'b0][1:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28, src/main/scala/snax/utils/Counter.scala:24:26[0J
      `endif // RANDOMIZE_REG_INIT[0J
      if (reset)	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
        value = 2'h0;	// src/main/scala/snax/utils/Counter.scala:24:26, :30:25[0J
    end // initial[0J
    `ifdef FIRRTL_AFTER_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.sca[0J[0Jla:100:28[0J
      `FIRRTL_AFTER_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28[0J
    `endif // FIRRTL_AFTER_INITIAL[0J
  `endif // ENABLE_INITIAL_REG_[0J
  assign io_value = value;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:28, src/main/scala/snax/utils/Counter.scala:24:26[0J
endmodule[0J
[0J
module RescaleDown_Anon(	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:25[0J
  input  [31:0] io_data_i_bits,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:12:14[0J
  output [7:0]  io_data_o,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:12:14[0J
  input  [31:0] io_input_zp,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:12:14[0J
                io_multiplier,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:12:14[0J
                io_output_zp,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:12:14[0J
  input  [7:0]  io_shift	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:12:14[0J
);[0J
[0J
  wire [31:0]  _zero_compensated_data_i_T = io_data_i_bits - io_input_zp;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:22:45[0J
  wire [256:0] _shifted_one_T_2 = 257'h1 << io_shift - 8'h1;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:28:{23,36}[0J
  wire [63:0]  _shifted_data_i_T =[0J
    {{32{_zero_compensated_data_i_T[31]}}, _zero_compensated_data_i_T}[0J
    * {32'h0, io_multiplier} + _shifted_one_T_2[63:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:22:45, :25:48, :28:{15,23}, :31:40[0J
  wire [63:0]  shifted_value =[0J
    $signed($signed((|(io_shift[7:5]))[0J
                      ? ($signed(_zero_compensated_data_i_T) > -32'sh1[0J
                           ? _shifted_data_i_T + 64'h40000000[0J
                           : _shifted_data_i_T - 64'h40000000)[0J
                      : _shifted_data_i_T) >>> io_shift);	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:22:45, :31:40, :34:{32,40}, :35:{20,38}, :37:{20,38}, :41:{17,25}, :42:25, :44:25, :48:40[0J
  wire [31:0]  _zero_compensated_out_T = shifted_value[31:0] + io_output_zp;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:48:40, :51:24, :54:48[0J
  assign io_data_o =[0J
    $signed(_zero_compensated_out_T) > 32'sh7F[0J
      ? 8'h7F[0J
      : $signed(_zero_compensated_out_T) < -32'sh80[0J
          ? 8'h80[0J
          : _zero_compensated_out_T[7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:54:48, :58:{29,74}, :59:21, :60:{35,80}, :61:21, :63:21, :124:25[0J
endmodule[0J
[0J
module unnamed_cluster_DataPathExtension_RescaleDown(	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
  input          clock,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
                 reset,	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
  input  [31:0]  io_csr_i_0,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
                 io_csr_i_1,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
                 io_csr_i_2,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
                 io_csr_i_3,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  input          io_start_i,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
                 io_bypass_i,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  output         io_data_i_ready,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  input          io_data_i_valid,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  input  [511:0] io_data_i_bits,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  input          io_data_o_ready,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  output         io_data_o_valid,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  output [511:0] io_data_o_bits,	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
  output         io_busy_o	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:52:14[0J
);[0J
[0J
  wire [7:0]   _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [7:0]   _PE_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
  wire [1:0]   _counter_io_value;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23[0J
  wire         _outputMux_io_in_1_ready;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:39[0J
  wire         _inputDemux_io_out_1_valid;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:40[0J
  wire [511:0] _inputDemux_io_out_1_bits;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:40[0J
  wire         ext_data_o_ready;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:66:24[0J
  wire         ext_data_i_ready = ext_data_o_ready;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, :66:24[0J
  wire         ext_data_i_valid;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24[0J
  wire         ext_busy_o;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:72:24[0J
  wire         _ext_data_o_valid_T = ext_data_i_ready & ext_data_i_valid;	// src/main/scala/chisel3/util/Decoupled.scala:51:35, src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24[0J
  assign ext_busy_o = |_counter_io_value;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:72:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :106:40[0J
  reg  [7:0]   regs_0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_1;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_2;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_3;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_4;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_5;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_6;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_7;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_8;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_9;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_10;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_11;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_12;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_13;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   reg[0J[0Js_14;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_15;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_16;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_17;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_18;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_19;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_20;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_21;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_22;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_23;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_24;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_25;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_26;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_27;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_28;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_29;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_30;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_31;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_32;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_33;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_34;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_35;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_36;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_37;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_38;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_39;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_40;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_41;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_42;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_43;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_44;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_45;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_46;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  reg  [7:0]   regs_47;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21[0J
  wire [511:0] ext_data_i_bits;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24[0J
  wire [511:0] ext_data_o_bits =[0J
    {_PE_15_io_data_o,[0J
     _PE_14_io_data_o,[0J
     _PE_13_io_data_o,[0J
     _PE_12_io_data_o,[0J
     _PE_11_io_data_o,[0J
     _PE_10_io_data_o,[0J
     _PE_9_io_data_o,[0J
     _PE_8_io_data_o,[0J
     _PE_7_io_data_o,[0J
     _PE_6_io_data_o,[0J
     _PE_5_io_data_o,[0J
     _PE_4_io_data_o,[0J
     _PE_3_io_data_o,[0J
     _PE_2_io_data_o,[0J
     _PE_1_io_data_o,[0J
     _PE_io_data_o,[0J
     regs_47,[0J
     regs_46,[0J
     regs_45,[0J
     regs_44,[0J
     regs_43,[0J
     regs_42,[0J
     regs_41,[0J
     regs_40,[0J
     regs_39,[0J
     regs_38,[0J
     regs_37,[0J
     regs_36,[0J
     regs_35,[0J
     regs_34,[0J
     regs_33,[0J
     regs_32,[0J
     regs_31,[0J
     regs_30,[0J
     regs_29,[0J
     regs_28,[0J
     regs_27,[0J
     regs_26,[0J
     regs_25,[0J
     regs_24,[0J
     regs_23,[0J
     regs_22,[0J
     regs_21,[0J
     regs_20,[0J
     regs_19,[0J
     regs_18,[0J
     regs_17,[0J
     regs_16,[0J
     regs_15,[0J
     regs_14,[0J
     regs_13,[0J
     regs_12,[0J
     regs_11,[0J
     regs_10,[0J
     regs_9,[0J
     regs_8,[0J
     regs_7,[0J
     regs_6,[0J
     regs_5,[0J
     regs_4,[0J
     regs_3,[0J
     regs_2,[0J
     regs_1,[0J
     regs_0};	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:66:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20, :147:58[0J
  wire         ext_data_o_valid = _ext_data_o_valid_T & (&_counter_io_value);	// src/main/scala/chisel3/util/Decoupled.scala:51:35, src/main/scala/snax/DataPathExtension/DataPathExtension.scala:66:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :148:{39,59}[0J
  always @(posedge clock or posedge reset) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
    if (reset) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
      regs_0 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_1 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_2 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_3 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_4 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_5 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_6 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_7 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_8 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_9 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_10 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_11 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_12 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_13 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_14 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_15 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_16 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_17 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_18 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_19 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_20 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_21 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_22 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_23 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_24 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_25 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_26 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_27 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_28 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_29 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_30 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_31 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_32 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_33 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_34 <= 8'h0;	// src/main/scala/s[0J[0Jnax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_35 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_36 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_37 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_38 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_39 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_40 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_41 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_42 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_43 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_44 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_45 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_46 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      regs_47 <= 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
    end[0J
    else if (_ext_data_o_valid_T) begin	// src/main/scala/chisel3/util/Decoupled.scala:51:35[0J
      automatic logic [5:0] _GEN = {_counter_io_value, 4'h0};	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :100:23, :141:80[0J
      automatic logic [5:0] _GEN_0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_1;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_2;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_3;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_4;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_5;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_6;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_7;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_8;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_9;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_10;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_11;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_12;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_13;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:80[0J
      automatic logic [5:0] _GEN_14 = _GEN + 6'hF;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_0 = _GEN + 6'h1;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_1 = _GEN + 6'h2;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_2 = _GEN + 6'h3;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_3 = _GEN + 6'h4;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_4 = _GEN + 6'h5;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_5 = _GEN + 6'h6;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_6 = _GEN + 6'h7;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_7 = _GEN + 6'h8;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_8 = _GEN + 6'h9;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_9 = _GEN + 6'hA;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_10 = _GEN + 6'hB;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_11 = _GEN + 6'hC;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_12 = _GEN + 6'hD;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      _GEN_13 = _GEN + 6'hE;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:141:{80,87}[0J
      if ((&_counter_io_value) | (|_GEN_14)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | (|_GEN_13)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | (|_GEN_12)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | (|_GEN_11)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | (|_GEN_10)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | (|_GEN_9)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | (|_GEN_8)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | (|_GEN_7)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | (|_GEN_6)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | (|_GEN_5)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | (|_GEN_4)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | (|_GEN_3)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | (|_GEN_2)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | (|_GEN_1)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | (|_GEN_0)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                    if ((&_counter_io_value) | (|_counter_io_value)) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :140:{29,81}, :141:87[0J
                                    end[0J
                                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :140:{29,81}, :141:87[0J
                                      regs_0 <= _PE_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_0 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_0 <= _PE_2_io_data_o;	// [0J[0Jsrc/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_0 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_0 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_0 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_0 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_0 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_0 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_0 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_0 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_0 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_0 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_0 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_0 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_0 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_1 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_1 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_1 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_1 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_1 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_1 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_1 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/sca[0J[0Jla/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_1 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_1 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_1 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_1 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_1 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_1 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_1 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_1 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_2 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_2 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_2 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_2 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_2 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_2 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_2 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_2 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_2 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_2 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_2 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_2 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_2 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
[0J          regs_2 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_2 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h3) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_3 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_3 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_3 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_3 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_3 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_3 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_3 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_3 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_3 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_3 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_3 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_3 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_3 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_3 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_3 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81},[0J[0J :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h4) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_4 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_4 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_4 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_4 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_4 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_4 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_4 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_4 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_4 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_4 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_4 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_4 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_4 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_4 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_4 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h5) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  [0J[0J                end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_5 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_5 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_5 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_5 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_5 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_5 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_5 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_5 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_5 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_5 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_5 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_5 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_5 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_5 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_5 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h6) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_6 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_6 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_6 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_6 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_6 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtens[0J[0Jion/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_6 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_6 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_6 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_6 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_6 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_6 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_6 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_6 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_6 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_6 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h7) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_7 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_7 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_7 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_7 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_7 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_7 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_7 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_7 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_7 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_7 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_7 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/[0J[0JRescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_7 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_7 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_7 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_7 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h8) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_8 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_8 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_8 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_8 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_8 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_8 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_8 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_8 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_8 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_8 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_8 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_8 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_8 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_8 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_8 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
      [0J[0J        if ((&_counter_io_value) | _GEN_10 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h9) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_9 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_9 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_9 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_9 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_9 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_9 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_9 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_9 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_9 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_9 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_9 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_9 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_9 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_9 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_9 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'hA) begin	// src[0J[0J/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'hA) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_10 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_10 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_10 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_10 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_10 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_10 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_10 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_10 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_10 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_10 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_10 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_10 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_10 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_10 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_10 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'hB) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_11 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_11 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_11 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27[0J[0J, :140:{29,81}, :141:87[0J
                              regs_11 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_11 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_11 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_11 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_11 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_11 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_11 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_11 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_11 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_11 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_11 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_11 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'hC) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_12 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_12 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_12 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_12 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_12 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_12 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_12 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_12 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_12 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J[0J[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_12 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_12 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_12 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_12 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_12 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_12 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'hD) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_13 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_13 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_13 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_13 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_13 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_13 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_13 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_13 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_13 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_13 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_13 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_13 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_13 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_13 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_13 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100[0J[0J:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'hE) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_14 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_14 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_14 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_14 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_14 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_14 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_14 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_14 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_14 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_14 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_14 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_14 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_14 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_14 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_14 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 ![0J[0J= 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'hF) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_15 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_15 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_15 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_15 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_15 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_15 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_15 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_15 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_15 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_15 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_15 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_15 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_15 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_15 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_15 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h10) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                    if ((&_counter_io_value)[0J
                                        | _counter_io_value != 2'h1) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :140:{29,81}, :141:87[0J
                                    end[0J
                                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :140:{29,81}, :141:87[0J
                     [0J[0J                 regs_16 <= _PE_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_16 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_16 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_16 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_16 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_16 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_16 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_16 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_16 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_16 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_16 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_16 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_16 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_16 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_16 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_16 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h11) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_17 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_17 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_17 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_17 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_17 <= _PE_5_io_data_o[0J[0J;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_17 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_17 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_17 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_17 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_17 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_17 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_17 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_17 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_17 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_17 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h12) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_18 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_18 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_18 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_18 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_18 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_18 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_18 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_18 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_18 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_18 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,[0J[0J81}, :141:87[0J
                regs_18 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_18 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_18 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_18 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_18 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h13) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_19 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_19 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_19 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_19 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_19 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_19 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_19 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_19 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_19 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_19 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_19 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_19 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_19 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_19 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_19 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/Rescale[0J[0JDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h14) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_20 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_20 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_20 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_20 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_20 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_20 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_20 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_20 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_20 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_20 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_20 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_20 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_20 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_20 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_20 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:[0J[0J{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h15) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_21 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_21 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_21 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_21 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_21 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_21 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_21 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_21 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_21 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_21 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_21 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_21 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_21 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_21 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_21 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h16) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_22 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_22 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.[0J[0Jscala:139:27, :140:{29,81}, :141:87[0J
                                regs_22 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_22 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_22 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_22 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_22 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_22 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_22 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_22 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_22 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_22 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_22 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_22 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_22 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h17) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_23 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_23 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_23 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_23 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_23 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_23 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_23 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_23 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExte[0J[0Jnsion/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_23 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_23 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_23 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_23 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_23 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_23 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_23 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h18) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_24 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_24 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_24 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_24 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_24 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_24 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_24 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_24 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_24 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_24 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_24 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_24 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_24 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_24 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J[0J[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_24 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h19) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_25 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_25 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_25 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_25 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_25 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_25 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_25 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_25 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_25 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_25 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_25 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_25 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_25 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_25 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_25 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1A) begin	[0J[0J// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_26 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_26 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_26 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_26 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_26 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_26 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_26 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_26 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_26 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_26 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_26 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_26 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_26 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_26 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_26 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                          [0J[0J        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_27 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_27 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_27 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_27 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_27 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_27 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_27 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_27 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_27 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_27 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_27 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_27 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_27 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_27 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_27 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_28 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_28 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_28 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_28 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_28 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/Rescale[0J[0JDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_28 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_28 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_28 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_28 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_28 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_28 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_28 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_28 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_28 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_28 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_29 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_29 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_29 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_29 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_29 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_29 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_29 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_29 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_29 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_29 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_29 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scal[0J[0Ja/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_29 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_29 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_29 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_29 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_30 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_30 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_30 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_30 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_30 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_30 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_30 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_30 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_30 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_30 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_30 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_30 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_30 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_30 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_30 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.sc[0J[0Jala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h1F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_31 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_31 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_31 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_31 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_31 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_31 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_31 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_31 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_31 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_31 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_31 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_31 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_31 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_31 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_31 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81[0J[0J}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h20) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                    if ((&_counter_io_value)[0J
                                        | _counter_io_value != 2'h2) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :140:{29,81}, :141:87[0J
                                    end[0J
                                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :140:{29,81}, :141:87[0J
                                      regs_32 <= _PE_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_32 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_32 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_32 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_32 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_32 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_32 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_32 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_32 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_32 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_32 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_32 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_32 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_32 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_32 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_32 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h21) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_33 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                        [0J[0J        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_33 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_33 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_33 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_33 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_33 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_33 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_33 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_33 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_33 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_33 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_33 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_33 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_33 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_33 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h22) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_34 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_34 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_34 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_34 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_34 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_34 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81[0J[0J}, :141:87[0J
                        regs_34 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_34 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_34 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_34 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_34 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_34 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_34 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_34 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_34 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h23) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_35 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_35 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_35 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_35 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_35 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_35 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_35 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_35 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_35 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_35 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_35 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_35 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, [0J[0J:141:87[0J
            regs_35 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_35 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_35 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h24) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_36 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_36 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_36 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_36 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_36 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_36 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_36 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_36 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_36 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_36 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_36 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_36 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_36 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_36 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_36 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h25) begin	/[0J[0J/ src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h25) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_37 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_37 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_37 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_37 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_37 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_37 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_37 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_37 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_37 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_37 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_37 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_37 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_37 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_37 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_37 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h26) begin	// src/main[0J[0J/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h26) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_38 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_38 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_38 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_38 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_38 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_38 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_38 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_38 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_38 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_38 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_38 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_38 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_38 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_38 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_38 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h27) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_39 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_39 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_39 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_39 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                         [0J[0J end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_39 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_39 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_39 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_39 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_39 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_39 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_39 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_39 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_39 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_39 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_39 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h28) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_40 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_40 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_40 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_40 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_40 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_40 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_40 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_40 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_40 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_40 <= _PE_10_io_data_o;	// src/ma[0J[0Jin/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_40 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_40 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_40 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_40 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_40 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h29) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_41 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_41 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_41 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_41 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_41 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_41 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_41 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_41 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_41 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_41 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_41 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_41 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_41 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_41 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_41 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/R[0J[0JescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2A) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_42 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_42 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_42 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_42 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_42 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_42 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_42 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_42 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_42 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_42 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_42 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_42 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_42 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_42 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_42 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
 [0J[0J                         if ((&_counter_io_value) | _GEN_4 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2B) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_43 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_43 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_43 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_43 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_43 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_43 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_43 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_43 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_43 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_43 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_43 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_43 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_43 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_43 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_43 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2C) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_44 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_44 <= _PE_2_io_data_o;	// src/main/scala/[0J[0Jsnax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_44 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_44 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_44 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_44 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_44 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_44 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_44 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_44 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_44 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_44 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_44 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_44 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_44 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2D) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_45 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_45 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_45 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_45 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_45 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_45 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_45 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    [0J[0Jelse	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_45 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_45 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_45 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_45 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_45 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_45 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_45 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_45 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2E) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_46 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_46 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_46 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_46 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_46 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_46 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_46 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_46 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_46 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_46 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_46 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_46 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_46 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathEx[0J[0Jtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_46 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_46 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      if ((&_counter_io_value) | _GEN_14 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
        if ((&_counter_io_value) | _GEN_13 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
          if ((&_counter_io_value) | _GEN_12 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
            if ((&_counter_io_value) | _GEN_11 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
              if ((&_counter_io_value) | _GEN_10 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                if ((&_counter_io_value) | _GEN_9 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                  if ((&_counter_io_value) | _GEN_8 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                    if ((&_counter_io_value) | _GEN_7 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                      if ((&_counter_io_value) | _GEN_6 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                        if ((&_counter_io_value) | _GEN_5 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                          if ((&_counter_io_value) | _GEN_4 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                            if ((&_counter_io_value) | _GEN_3 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                              if ((&_counter_io_value) | _GEN_2 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                if ((&_counter_io_value) | _GEN_1 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  if ((&_counter_io_value) | _GEN_0 != 6'h2F) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23, :113:21, :139:27, :140:{29,81}, :141:{80,87}[0J
                                  end[0J
                                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                    regs_47 <= _PE_1_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                                end[0J
                                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                  regs_47 <= _PE_2_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                              end[0J
                              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                                regs_47 <= _PE_3_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                            end[0J
                            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                              regs_47 <= _PE_4_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                          end[0J
                          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                            regs_47 <= _PE_5_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                        end[0J
                        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                          regs_47 <= _PE_6_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                      end[0J
                      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                        regs_47 <= _PE_7_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                    end[0J
                    else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                      regs_47 <= _PE_8_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                  end[0J
                  else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                    regs_47 <= _PE_9_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
                end[0J
                else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                  regs_47 <= _PE_10_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
              end[0J
              else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
                regs_47 <= _PE_11_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
            end[0J
            else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
              regs_47 <= _PE_12_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
          end[0J
          else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
            regs_47 <= _PE_13_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
        end[0J
        else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
          regs_47 <= _PE_14_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
      end[0J
      else	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:139:27, :140:{29,81}, :141:87[0J
        regs_47 <= _PE_15_io_data_o;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :124:20[0J
    end[0J
  end // always @(posedge, posedge)[0J
  `ifdef ENABLE_INITIAL_REG_	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
    `ifdef FIRRTL_BEFORE_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
      `FIRRTL_BEFORE_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
    `endif // FIRRTL_BEFORE_INITIAL[0J
    initial begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
      automatic logic [31:0] _RANDOM[0:11];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
      `ifdef INIT_RANDOM_PROLOG_	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
        `INIT_RANDOM_PROLOG_	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
      `endif // INIT_RANDOM_PROLOG_[0J
      `ifdef RANDOMIZE_REG_INIT	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
        for (logic [3:0] i = 4'h0; i < 4'hC; i += 4'h1) begin[0J
          _RANDOM[i] = `RANDOM;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
        end	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:7[0J[0J8:11[0J
        regs_0 = _RANDOM[4'h0][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_1 = _RANDOM[4'h0][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_2 = _RANDOM[4'h0][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_3 = _RANDOM[4'h0][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_4 = _RANDOM[4'h1][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_5 = _RANDOM[4'h1][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_6 = _RANDOM[4'h1][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_7 = _RANDOM[4'h1][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_8 = _RANDOM[4'h2][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_9 = _RANDOM[4'h2][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_10 = _RANDOM[4'h2][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_11 = _RANDOM[4'h2][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_12 = _RANDOM[4'h3][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_13 = _RANDOM[4'h3][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_14 = _RANDOM[4'h3][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_15 = _RANDOM[4'h3][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_16 = _RANDOM[4'h4][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_17 = _RANDOM[4'h4][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_18 = _RANDOM[4'h4][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_19 = _RANDOM[4'h4][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_20 = _RANDOM[4'h5][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_21 = _RANDOM[4'h5][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_22 = _RANDOM[4'h5][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_23 = _RANDOM[4'h5][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_24 = _RANDOM[4'h6][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_25 = _RANDOM[4'h6][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_26 = _RANDOM[4'h6][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_27 = _RANDOM[4'h6][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_28 = _RANDOM[4'h7][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_29 = _RANDOM[4'h7][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_30 = _RANDOM[4'h7][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_31 = _RANDOM[4'h7][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_32 = _RANDOM[4'h8][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_33 = _RANDOM[4'h8][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_34 = _RANDOM[4'h8][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_35 = _RANDOM[4'h8][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_36 = _RANDOM[4'h9][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_37 = _RANDOM[4'h9][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_38 = _RANDOM[4'h9][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_39 = _RANDOM[4'h9][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_40 = _RANDOM[4'hA][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_41 = _RANDOM[4'hA][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_42 = _RANDOM[4'hA][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_43 = _RANDOM[4'hA][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_44 = _RANDOM[4'hB][7:0];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_45 = _RANDOM[4'hB][15:8];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_46 = _RANDOM[4'hB][23:16];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
        regs_47 = _RANDOM[4'hB][31:24];	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11, :113:21[0J
      `endif // RANDOMIZE_REG_INIT[0J
      if (reset) begin	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
        regs_0 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_1 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_2 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_3 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_4 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_5 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_6 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_7 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_8 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_9 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_10 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_11 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_12 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_13 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_14 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_15 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_16 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_17 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_18 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_19 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_20 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_21 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_22 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_23 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_24 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_25 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_26 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDo[0J[0Jwn.scala:113:21, :114:12[0J
        regs_27 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_28 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_29 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_30 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_31 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_32 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_33 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_34 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_35 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_36 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_37 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_38 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_39 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_40 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_41 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_42 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_43 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_44 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_45 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_46 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
        regs_47 = 8'h0;	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:113:21, :114:12[0J
      end[0J
    end // initial[0J
    `ifdef FIRRTL_AFTER_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
      `FIRRTL_AFTER_INITIAL	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
    `endif // FIRRTL_AFTER_INITIAL[0J
  `endif // ENABLE_INITIAL_REG_[0J
  DataPathExtension_Demux_W512 inputDemux (	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:40[0J
    .io_in_ready    (io_data_i_ready),[0J
    .io_in_valid    (io_data_i_valid),[0J
    .io_in_bits     (io_data_i_bits),[0J
    .io_out_0_ready (ext_data_i_ready),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24[0J
    .io_out_0_valid (ext_data_i_valid),[0J
    .io_out_0_bits  (ext_data_i_bits),[0J
    .io_out_1_ready (_outputMux_io_in_1_ready),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:39[0J
    .io_out_1_valid (_inputDemux_io_out_1_valid),[0J
    .io_out_1_bits  (_inputDemux_io_out_1_bits),[0J
    .io_sel         (io_bypass_i)[0J
  );[0J
  DataPathExtension_Mux_W512 outputMux (	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:88:39[0J
    .io_in_0_ready (ext_data_o_ready),[0J
    .io_in_0_valid (ext_data_o_valid),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:66:24[0J
    .io_in_0_bits  (ext_data_o_bits),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:66:24[0J
    .io_in_1_ready (_outputMux_io_in_1_ready),[0J
    .io_in_1_valid (_inputDemux_io_out_1_valid),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:40[0J
    .io_in_1_bits  (_inputDemux_io_out_1_bits),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:77:40[0J
    .io_out_ready  (io_data_o_ready),[0J
    .io_out_valid  (io_data_o_valid),[0J
    .io_out_bits   (io_data_o_bits),[0J
    .io_sel        (io_bypass_i)[0J
  );[0J
  RescaleDownCounter counter (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:100:23[0J
    .clock    (clock),[0J
    .reset    (reset),[0J
    .io_tick  (_ext_data_o_valid_T),	// src/main/scala/chisel3/util/Decoupled.scala:51:35[0J
    .io_reset (io_start_i),[0J
    .io_value (_counter_io_value)[0J
  );[0J
  RescaleDown_Anon PE (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[31:0]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_1 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[63:32]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_1_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_2 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[95:64]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_2_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_3 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[127:96]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_3_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_4 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[159:128]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_4_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_5 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[191:160]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_5_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_6 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[223:192]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_6_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_7 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[255:224]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_7_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .i[0J[0Jo_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_8 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[287:256]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_8_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_9 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[319:288]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_9_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_10 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[351:320]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_10_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_11 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[383:352]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_11_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_12 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[415:384]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_12_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_13 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[447:416]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_13_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_14 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[479:448]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_14_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  RescaleDown_Anon PE_15 (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:124:20[0J
    .io_data_i_bits (ext_data_i_bits[511:480]),	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, src/main/scala/snax/DataPathExtension/RescaleDown.scala:129:12[0J
    .io_data_o      (_PE_15_io_data_o),[0J
    .io_input_zp    (io_csr_i_0),[0J
    .io_multiplier  (io_csr_i_1),[0J
    .io_output_zp   (io_csr_i_2),[0J
    .io_shift       (io_csr_i_3[7:0])	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:137:24[0J
  );[0J
  assign io_busy_o = ext_busy_o | ext_data_i_valid;	// src/main/scala/snax/DataPathExtension/DataPathExtension.scala:64:24, :72:24, :74:27, src/main/scala/snax/DataPathExtension/RescaleDown.scala:78:11[0J
endmodule[0J
[0J
module unnamed_cluster_DataPathExtensionHost(	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:37:7[0J
  input          clock,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:37:7[0J
                 reset,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:37:7[0J
  output         io_data_in_ready,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  input          io_data_in_valid,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  input  [511:0] io_data_in_bits,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  input          io_data_out_ready,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  output         io_data_out_valid,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  output [511:0] io_data_out_bits,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  input          io_cfg_bypass,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  input  [31:0]  io_cfg_userCsr_0,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
                 io_cfg_userCsr_1,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
                 io_cfg_userCsr_2,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
                 io_cfg_userCsr_3,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  input          io_start,	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
  output         io_busy	// src/main/scala/snax/DataPathExtension/DataPathExtensionHost.scala:46:32[0J
);[0J
[0J
  unnamed_cluster_DataPathExtension_RescaleDown unnamed_cluster_Extension_0_RescaleDown (	// src/main/scala/snax/DataPathExtension/RescaleDown.scala:77:11[0J
    .clock           (clock),[0J
    .reset           (reset),[0J
    .io_csr_i_0      (io_cfg_userCsr_0),[0J
    .io_csr_i_1      (io_cfg_userCsr_1),[0J
    .io_csr_i_2      (io_cfg_userCsr_2),[0J
    .io_csr_i_3      (io_cfg_userCsr_3),[0J
    .io_start_i      (io_start),[0J
    .io_bypass_i     (io_cfg_bypass),[0J
    .io_data_i_ready (io_data_in_ready),[0J
    .io_data_i_valid (io_data_in_valid),[0J
    .io_data_i_bits  (io_data_in_bits),[0J
    .io_data_o_ready (io_data_out_ready),[0J
    .io_data_o_valid (io_data_out_valid),[0J
    .io_data_o_bits  (io_data_out_bits),[0J
    .io_busy_o       (io_busy)[0J
  );[0J
endmodule[0J
[0J
[0J[0J[0J[0m[[0m[32msuccess[0m] [0m[0mTotal time: 10 s, completed Aug 4, 2025, 3:01:16 PM[0m[0J
[0J[0J